`timescale 1ms/10ps
module tb;


endmodule