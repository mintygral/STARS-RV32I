`timescale 1ms/10ps

module tb_register_file;

endmodule